`include "test_with_port.sv"
`include "design.sv"
`include "top.sv"