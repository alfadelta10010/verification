module test;
real r5;
shortreal r6;
initial
begin
r5 = 6.777;
r6 = 3.1;
$display(r5, " ", r6);
end
endmodule