`include "test_with_mp.sv"
`include "design.sv"
`include "top.sv"
`include "ifc.sv"